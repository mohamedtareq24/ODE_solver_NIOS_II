module memo_interface (
    input read ,input  [8:0] Data_in ,
    output reg [8:0] Data_out 
);
VGA_interface Controller()
register  Memory()
endmodule //memo_interface